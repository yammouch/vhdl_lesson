library ieee;
use ieee.std_logic_1164.all;

entity sub1 is
  port (
    pulse : in std_ulogic );
end entity;
