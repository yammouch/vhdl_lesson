library ieee;
use ieee.std_logic_1164.all;

entity sim_top is
end entity;

architecture sim1 of sim_top is
begin
  process
  begin
    report "sim1";
    wait;
  end process;
end sim1;
